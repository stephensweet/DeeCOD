
/* 
 not gate
*/
module gatedesign
(
 a,
 out
 );

   input a;

   output out;

 assign out = ~a;
 
endmodule // not_gate
